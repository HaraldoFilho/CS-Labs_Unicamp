Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;

entity tb_ALU is
end tb_ALU;

architecture behav of tb_ALU is

Component ALU is
	port(SrcA 	: in std_logic_vector(31 downto 0);
		SrcB 	: in std_logic_vector(31 downto 0);
		AluControl: in std_logic_vector(3 downto 0);
		AluResult : out std_logic_vector(31 downto 0);
		Zero 	: out std_logic;
		Overflow 	: out std_logic);
End Component;

for ALU_TB: ALU use entity work.ALU;
signal SrcA 		: std_logic_vector(31 downto 0);
signal SrcB 		: std_logic_vector(31 downto 0);
signal AluControl 	: std_logic_vector(3 downto 0);
signal AluResult 	: std_logic_vector(31 downto 0);
signal Zero 		: std_logic;
signal Overflow 	: std_logic;
 
Begin
	ALU_TB : ALU port map (SrcA, SrcB, AluControl, AluResult, Zero, Overflow);

	AluControl <= "0000", 			 
			    "0001" after 80 ns,    
			    "0010" after 160 ns,    
			    "0011" after 240 ns,   
			    "0100" after 320 ns,   
			    "0101" after 360 ns,   
			    "0110" after 400 ns,  
			    "0111" after 440 ns,
			    "1010" after 480 ns,   
			    "1011" after 540 ns,
			    "1111" after 600 ns;
	
	SrcA <= "00000000000000000000000000000000",
		   "11111111111111111111111111111111" after 20 ns,
		   "01111111111111111111111111111111" after 40 ns,
		   "00111110000000111111000000111110" after 60 ns,
		   "00000000000000000000000000000000" after 80 ns,
		   "11111111111111111111111111111111" after 100 ns,
		   "01111111111111111111111111111111" after 120 ns,
		   "00111110000000111111000000111110" after 140 ns,

		   "00000000000000000000000000000000" after 160 ns,
		   "11111111111111111111111111111111" after 180 ns,
		   "01111111111111111111111111111111" after 200 ns,
		   "00111110000000111111000000111110" after 220 ns,
		   "00000000000000000000000000000000" after 240 ns,
		   "11111111111111111111111111111111" after 260 ns,
		   "01111111111111111111111111111111" after 280 ns,
		   "00111110000000111111000000111110" after 300 ns,
	
		   "00000000000000000000000000000000" after 320 ns,
		   "11111111111111111111111111111111" after 330 ns,
	   	   "00000000000000000000000000000000" after 340 ns,
	   	   "11111111111111111111111111111111" after 350 ns,
		   "00000000000000000000000000000000" after 360 ns,
		   "11111111111111111111111111111111" after 370 ns,
	   	   "00000000000000000000000000000000" after 380 ns,
	   	   "11111111111111111111111111111111" after 390 ns,
		   "00000000000000000000000000000000" after 400 ns,
		   "11111111111111111111111111111111" after 410 ns,
	   	   "00000000000000000000000000000000" after 420 ns,
	   	   "11111111111111111111111111111111" after 430 ns,
		   "00000000000000000000000000000000" after 440 ns,
		   "11111111111111111111111111111111" after 450 ns,
	   	   "00000000000000000000000000000000" after 460 ns,
	   	   "11111111111111111111111111111111" after 470 ns,
		   "00000000000000000000000000000001" after 480 ns,
		   "00000000000000000000000000000010" after 490 ns,
		   "00000000000000000000000000000000" after 500 ns,
		   "11111111111111111111111111111111" after 510 ns,
		   "00000000000000000000000000000000" after 520 ns,
		   "11111111111111111111111111111111" after 530 ns,	
		   "00000000000000000000000000000001" after 540 ns,
		   "00000000000000000000000000000010" after 550 ns,
		   "00000000000000000000000000000000" after 560 ns,
		   "11111111111111111111111111111111" after 570 ns,
		   "00000000000000000000000000000000" after 580 ns,
		   "11111111111111111111111111111111" after 590 ns;	
		   
	SrcB <= "00000000000000000000000000000000" ,
		   "10000000000000000000000000000000" after 10 ns,
		   "11111111111111111111111111111111" after 20 ns,
		   "00000000000000000000000000000000" after 30 ns,
		   "00000000000000000000000000000001" after 40 ns,
		   "00000000000000000000000000000000" after 50 ns,
		   "11111100000111100000011100000111" after 60 ns,
		   "00000000000000000000000000000000" after 80 ns,
		   "10000000000000000000000000000000" after 90 ns,
		   "11111111111111111111111111111111" after 100 ns,
		   "00000000000000000000000000000000" after 110 ns,
		   "00000000000000000000000000000001" after 120 ns,
		   "00000000000000000000000000000000" after 130 ns,
		   "11111100000111100000011100000111" after 140 ns,

		   "00000000000000000000000000000000" after 160 ns,
		   "10000000000000000000000000000000" after 170 ns,
		   "11111111111111111111111111111111" after 180 ns,
		   "00000000000000000000000000000000" after 190 ns,
		   "00000000000000000000000000000001" after 200 ns,
		   "00000000000000000000000000000000" after 210 ns,
		   "11111100000111100000011100000111" after 220 ns,
		   "00000000000000000000000000000000" after 240 ns,
		   "10000000000000000000000000000000" after 250 ns,
		   "11111111111111111111111111111111" after 260 ns,
		   "00000000000000000000000000000000" after 270 ns,
		   "00000000000000000000000000000001" after 280 ns,
		   "00000000000000000000000000000000" after 290 ns,
		   "11111100000111100000011100000111" after 300 ns,
		   
		   "00000000000000000000000000000000" after 320 ns,	
		   "11111111111111111111111111111111" after 340 ns,
		   "00000000000000000000000000000000" after 360 ns,	
		   "11111111111111111111111111111111" after 380 ns,
		   "00000000000000000000000000000000" after 400 ns,	
		   "11111111111111111111111111111111" after 420 ns,
		   "00000000000000000000000000000000" after 440 ns,	
		   "11111111111111111111111111111111" after 460 ns,
		   "00000000000000000000000000000010" after 480 ns,
		   "00000000000000000000000000000001" after 500 ns,
		   "11111111111111111111111111111111" after 520 ns,
		   "00000000000000000000000000000010" after 540 ns,
		   "00000000000000000000000000000001" after 560 ns,
		   "11111111111111111111111111111111" after 580 ns;

End  behav;
